//==============================================================================
// QEDMMA IMM (Interacting Multiple Model) Tracker
// Author: Dr. Mladen Mešter
// Copyright (c) 2026 Dr. Mladen Mešter - All Rights Reserved
//
// Description:
//   Implements IMM filter with 3 motion models for robust target tracking:
//   - CV (Constant Velocity)
//   - CA (Constant Acceleration)  
//   - CT (Coordinated Turn)
//
//   - 9-state tracking (position, velocity, acceleration)
//   - Model probability adaptation
//   - Covariance intersection for track fusion
//   - FPGA-optimized fixed-point arithmetic
//
// References:
//   - [REQ-TRK-001] Track 50+ simultaneous targets
//   - [REQ-TRK-002] Maneuvering target tracking (up to 9g)
//   - [REQ-TRK-003] Track update rate ≥ 10 Hz
//
// Author: Dr. Mladen Mešter / Forge Swarm
// Date: 2026-01-31
// Version: 1.0
//==============================================================================

`timescale 1ns / 1ps

module imm_tracker #(
    // State vector parameters
    parameter int STATE_WIDTH    = 32,       // State component width
    parameter int FRAC_BITS      = 16,       // Fixed-point fractional bits
    parameter int MEAS_WIDTH     = 32,       // Measurement width
    
    // Filter parameters
    parameter int NUM_MODELS     = 3,        // Number of motion models
    parameter int STATE_DIM      = 9,        // State dimension [x,y,z,vx,vy,vz,ax,ay,az]
    parameter int MEAS_DIM       = 3,        // Measurement dimension [x,y,z]
    
    // Track management
    parameter int MAX_TRACKS     = 64,       // Maximum simultaneous tracks
    parameter int TRACK_ID_WIDTH = 8         // Track ID width
)(
    // Clock and reset
    input  logic                        clk,
    input  logic                        rst_n,
    
    // Measurement input
    input  logic [MEAS_DIM-1:0][MEAS_WIDTH-1:0] measurement,
    input  logic [15:0]                         meas_variance,   // Measurement noise
    input  logic                                meas_valid,
    
    // Track association input (from correlator)
    input  logic [TRACK_ID_WIDTH-1:0]           assoc_track_id,
    input  logic                                assoc_valid,
    input  logic                                new_track,       // Create new track
    
    // State output (selected track)
    output logic [STATE_DIM-1:0][STATE_WIDTH-1:0] state_out,
    output logic [STATE_DIM-1:0][STATE_WIDTH-1:0] covariance_diag, // Diagonal only
    output logic [TRACK_ID_WIDTH-1:0]             track_id_out,
    output logic                                  track_valid,
    
    // Model probabilities output
    output logic [NUM_MODELS-1:0][15:0]           model_probs,    // Fixed-point [0,1]
    
    // Track management output
    output logic [5:0]                            num_active_tracks,
    output logic                                  track_lost,
    output logic                                  track_confirmed,
    
    // Configuration
    input  logic [15:0]                           cfg_process_noise,
    input  logic [15:0]                           cfg_gate_threshold,
    input  logic [7:0]                            cfg_confirm_hits,
    input  logic [7:0]                            cfg_delete_misses,
    
    // Status
    output logic                                  busy,
    output logic                                  overflow
);

    //--------------------------------------------------------------------------
    // Model transition probability matrix (fixed)
    // π[i][j] = P(model j at k | model i at k-1)
    //--------------------------------------------------------------------------
    // Typical values: stay in same model with high probability
    localparam logic [15:0] PI_STAY  = 16'hCCCC;  // 0.8 in Q0.16
    localparam logic [15:0] PI_TRANS = 16'h1999;  // 0.1 in Q0.16
    
    //--------------------------------------------------------------------------
    // State machine
    //--------------------------------------------------------------------------
    typedef enum logic [3:0] {
        ST_IDLE,
        ST_RECEIVE_MEAS,
        ST_MIXING,
        ST_PREDICT_CV,
        ST_PREDICT_CA,
        ST_PREDICT_CT,
        ST_UPDATE_CV,
        ST_UPDATE_CA,
        ST_UPDATE_CT,
        ST_COMBINE,
        ST_TRACK_MGMT,
        ST_OUTPUT
    } state_t;
    
    state_t state, next_state;
    
    //--------------------------------------------------------------------------
    // Track memory (BRAM-based in real implementation)
    //--------------------------------------------------------------------------
    // Per-track state for each model
    typedef struct packed {
        logic [STATE_DIM-1:0][STATE_WIDTH-1:0] state;
        logic [STATE_DIM-1:0][STATE_WIDTH-1:0] covariance;  // Diagonal
        logic [15:0] probability;  // Model probability
    } model_state_t;
    
    typedef struct packed {
        logic                      active;
        logic [7:0]                hit_count;
        logic [7:0]                miss_count;
        logic                      confirmed;
        model_state_t              models [NUM_MODELS-1:0];
        logic [STATE_WIDTH-1:0]    combined_state [STATE_DIM-1:0];
    } track_t;
    
    track_t tracks [0:MAX_TRACKS-1];
    
    // Current working track
    logic [TRACK_ID_WIDTH-1:0] current_track_id;
    track_t current_track;
    
    //--------------------------------------------------------------------------
    // Model-specific process noise covariance
    //--------------------------------------------------------------------------
    logic [STATE_WIDTH-1:0] Q_cv [0:STATE_DIM-1];   // CV process noise
    logic [STATE_WIDTH-1:0] Q_ca [0:STATE_DIM-1];   // CA process noise  
    logic [STATE_WIDTH-1:0] Q_ct [0:STATE_DIM-1];   // CT process noise
    
    // Initialize process noise (scaled by cfg_process_noise)
    always_ff @(posedge clk) begin
        // CV: Low acceleration noise
        Q_cv[0] <= cfg_process_noise << 4;   // Position
        Q_cv[1] <= cfg_process_noise << 4;
        Q_cv[2] <= cfg_process_noise << 4;
        Q_cv[3] <= cfg_process_noise << 8;   // Velocity
        Q_cv[4] <= cfg_process_noise << 8;
        Q_cv[5] <= cfg_process_noise << 8;
        Q_cv[6] <= cfg_process_noise;        // Acceleration (low for CV)
        Q_cv[7] <= cfg_process_noise;
        Q_cv[8] <= cfg_process_noise;
        
        // CA: Medium acceleration noise
        Q_ca[0] <= cfg_process_noise << 4;
        Q_ca[1] <= cfg_process_noise << 4;
        Q_ca[2] <= cfg_process_noise << 4;
        Q_ca[3] <= cfg_process_noise << 6;
        Q_ca[4] <= cfg_process_noise << 6;
        Q_ca[5] <= cfg_process_noise << 6;
        Q_ca[6] <= cfg_process_noise << 10;  // High for CA
        Q_ca[7] <= cfg_process_noise << 10;
        Q_ca[8] <= cfg_process_noise << 10;
        
        // CT: High lateral acceleration noise
        Q_ct[0] <= cfg_process_noise << 4;
        Q_ct[1] <= cfg_process_noise << 4;
        Q_ct[2] <= cfg_process_noise << 4;
        Q_ct[3] <= cfg_process_noise << 8;
        Q_ct[4] <= cfg_process_noise << 8;
        Q_ct[5] <= cfg_process_noise << 6;   // Lower vertical
        Q_ct[6] <= cfg_process_noise << 12;  // Very high lateral
        Q_ct[7] <= cfg_process_noise << 12;
        Q_ct[8] <= cfg_process_noise << 8;
    end
    
    //--------------------------------------------------------------------------
    // State Machine
    //--------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= ST_IDLE;
        end else begin
            state <= next_state;
        end
    end
    
    always_comb begin
        next_state = state;
        
        case (state)
            ST_IDLE: begin
                if (meas_valid && assoc_valid) begin
                    next_state = ST_RECEIVE_MEAS;
                end
            end
            
            ST_RECEIVE_MEAS: begin
                next_state = ST_MIXING;
            end
            
            ST_MIXING: begin
                next_state = ST_PREDICT_CV;
            end
            
            ST_PREDICT_CV: begin
                next_state = ST_PREDICT_CA;
            end
            
            ST_PREDICT_CA: begin
                next_state = ST_PREDICT_CT;
            end
            
            ST_PREDICT_CT: begin
                next_state = ST_UPDATE_CV;
            end
            
            ST_UPDATE_CV: begin
                next_state = ST_UPDATE_CA;
            end
            
            ST_UPDATE_CA: begin
                next_state = ST_UPDATE_CT;
            end
            
            ST_UPDATE_CT: begin
                next_state = ST_COMBINE;
            end
            
            ST_COMBINE: begin
                next_state = ST_TRACK_MGMT;
            end
            
            ST_TRACK_MGMT: begin
                next_state = ST_OUTPUT;
            end
            
            ST_OUTPUT: begin
                next_state = ST_IDLE;
            end
            
            default: next_state = ST_IDLE;
        endcase
    end
    
    //--------------------------------------------------------------------------
    // Measurement Latching
    //--------------------------------------------------------------------------
    logic [MEAS_DIM-1:0][MEAS_WIDTH-1:0] meas_latched;
    logic [15:0] meas_var_latched;
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            meas_latched <= '0;
            meas_var_latched <= '0;
            current_track_id <= '0;
        end else if (state == ST_RECEIVE_MEAS) begin
            meas_latched <= measurement;
            meas_var_latched <= meas_variance;
            current_track_id <= assoc_track_id;
            
            if (new_track) begin
                // Initialize new track
                current_track.active <= 1'b1;
                current_track.hit_count <= 8'd1;
                current_track.miss_count <= 8'd0;
                current_track.confirmed <= 1'b0;
                
                // Initialize all models with measurement
                for (int m = 0; m < NUM_MODELS; m++) begin
                    current_track.models[m].state[0] <= measurement[0];
                    current_track.models[m].state[1] <= measurement[1];
                    current_track.models[m].state[2] <= measurement[2];
                    for (int i = 3; i < STATE_DIM; i++) begin
                        current_track.models[m].state[i] <= '0;
                    end
                    current_track.models[m].probability <= 16'h5555;  // 1/3
                end
            end else begin
                current_track <= tracks[assoc_track_id];
            end
        end
    end
    
    //--------------------------------------------------------------------------
    // IMM Mixing Step
    // Mixed state: x̄_j = Σ_i μ_{i|j} * x̂_i
    // where μ_{i|j} = (1/c_j) * π_{ij} * μ_i
    //--------------------------------------------------------------------------
    logic [STATE_DIM-1:0][STATE_WIDTH-1:0] mixed_states [NUM_MODELS-1:0];
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int m = 0; m < NUM_MODELS; m++) begin
                for (int i = 0; i < STATE_DIM; i++) begin
                    mixed_states[m][i] <= '0;
                end
            end
        end else if (state == ST_MIXING) begin
            // Simplified mixing: weighted average based on transition probabilities
            for (int j = 0; j < NUM_MODELS; j++) begin
                for (int s = 0; s < STATE_DIM; s++) begin
                    automatic logic signed [2*STATE_WIDTH-1:0] sum = '0;
                    for (int i = 0; i < NUM_MODELS; i++) begin
                        // μ_{i|j} * x̂_i (simplified using stay/trans probabilities)
                        if (i == j) begin
                            sum = sum + ($signed(current_track.models[i].state[s]) * 
                                        $signed({16'b0, PI_STAY}));
                        end else begin
                            sum = sum + ($signed(current_track.models[i].state[s]) * 
                                        $signed({16'b0, PI_TRANS}));
                        end
                    end
                    mixed_states[j][s] <= sum[STATE_WIDTH+15:16];  // Normalize
                end
            end
        end
    end
    
    //--------------------------------------------------------------------------
    // Kalman Prediction (per model)
    // x̄ = F * x
    // P̄ = F * P * F' + Q
    //--------------------------------------------------------------------------
    logic [STATE_DIM-1:0][STATE_WIDTH-1:0] predicted_states [NUM_MODELS-1:0];
    logic [STATE_DIM-1:0][STATE_WIDTH-1:0] predicted_cov [NUM_MODELS-1:0];
    
    // Time step (100 ms = 0.1s, represented in fixed-point)
    localparam logic [STATE_WIDTH-1:0] DT = 32'h00001999;  // 0.1 in Q16.16
    
    // CV Prediction: x(k+1) = x(k) + v*dt, v(k+1) = v(k)
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int i = 0; i < STATE_DIM; i++) begin
                predicted_states[0][i] <= '0;
                predicted_cov[0][i] <= '0;
            end
        end else if (state == ST_PREDICT_CV) begin
            // Position: x += v * dt
            predicted_states[0][0] <= mixed_states[0][0] + 
                ((mixed_states[0][3] * DT) >>> FRAC_BITS);
            predicted_states[0][1] <= mixed_states[0][1] + 
                ((mixed_states[0][4] * DT) >>> FRAC_BITS);
            predicted_states[0][2] <= mixed_states[0][2] + 
                ((mixed_states[0][5] * DT) >>> FRAC_BITS);
            
            // Velocity: constant
            predicted_states[0][3] <= mixed_states[0][3];
            predicted_states[0][4] <= mixed_states[0][4];
            predicted_states[0][5] <= mixed_states[0][5];
            
            // Acceleration: zero for CV
            predicted_states[0][6] <= '0;
            predicted_states[0][7] <= '0;
            predicted_states[0][8] <= '0;
            
            // Covariance prediction (simplified diagonal update)
            for (int i = 0; i < STATE_DIM; i++) begin
                predicted_cov[0][i] <= current_track.models[0].covariance[i] + Q_cv[i];
            end
        end
    end
    
    // CA Prediction: x += v*dt + 0.5*a*dt^2, v += a*dt, a = const
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int i = 0; i < STATE_DIM; i++) begin
                predicted_states[1][i] <= '0;
                predicted_cov[1][i] <= '0;
            end
        end else if (state == ST_PREDICT_CA) begin
            // Position: x += v*dt + 0.5*a*dt^2
            logic signed [2*STATE_WIDTH-1:0] dt_sq;
            dt_sq = (DT * DT) >>> FRAC_BITS;
            
            predicted_states[1][0] <= mixed_states[1][0] + 
                ((mixed_states[1][3] * DT) >>> FRAC_BITS) +
                ((mixed_states[1][6] * dt_sq) >>> (FRAC_BITS + 1));
            predicted_states[1][1] <= mixed_states[1][1] + 
                ((mixed_states[1][4] * DT) >>> FRAC_BITS) +
                ((mixed_states[1][7] * dt_sq) >>> (FRAC_BITS + 1));
            predicted_states[1][2] <= mixed_states[1][2] + 
                ((mixed_states[1][5] * DT) >>> FRAC_BITS) +
                ((mixed_states[1][8] * dt_sq) >>> (FRAC_BITS + 1));
            
            // Velocity: v += a*dt
            predicted_states[1][3] <= mixed_states[1][3] + 
                ((mixed_states[1][6] * DT) >>> FRAC_BITS);
            predicted_states[1][4] <= mixed_states[1][4] + 
                ((mixed_states[1][7] * DT) >>> FRAC_BITS);
            predicted_states[1][5] <= mixed_states[1][5] + 
                ((mixed_states[1][8] * DT) >>> FRAC_BITS);
            
            // Acceleration: constant
            predicted_states[1][6] <= mixed_states[1][6];
            predicted_states[1][7] <= mixed_states[1][7];
            predicted_states[1][8] <= mixed_states[1][8];
            
            // Covariance
            for (int i = 0; i < STATE_DIM; i++) begin
                predicted_cov[1][i] <= current_track.models[1].covariance[i] + Q_ca[i];
            end
        end
    end
    
    // CT Prediction (simplified - real CT uses turn rate state)
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int i = 0; i < STATE_DIM; i++) begin
                predicted_states[2][i] <= '0;
                predicted_cov[2][i] <= '0;
            end
        end else if (state == ST_PREDICT_CT) begin
            // Similar to CA but with higher lateral uncertainty
            predicted_states[2] <= predicted_states[1];  // Use CA prediction
            
            // Higher covariance for maneuvering
            for (int i = 0; i < STATE_DIM; i++) begin
                predicted_cov[2][i] <= current_track.models[2].covariance[i] + Q_ct[i];
            end
        end
    end
    
    //--------------------------------------------------------------------------
    // Kalman Update (per model)
    // Innovation: y = z - H*x̄
    // Kalman gain: K = P̄*H' / (H*P̄*H' + R)
    // Updated state: x = x̄ + K*y
    // Updated covariance: P = (I - K*H)*P̄
    //--------------------------------------------------------------------------
    logic [STATE_DIM-1:0][STATE_WIDTH-1:0] updated_states [NUM_MODELS-1:0];
    logic [STATE_DIM-1:0][STATE_WIDTH-1:0] updated_cov [NUM_MODELS-1:0];
    logic [NUM_MODELS-1:0][31:0] likelihoods;
    
    // Update for each model (CV, CA, CT have same measurement model H = [I 0 0])
    genvar m;
    generate
        for (m = 0; m < NUM_MODELS; m++) begin : gen_update
            always_ff @(posedge clk or negedge rst_n) begin
                if (!rst_n) begin
                    for (int i = 0; i < STATE_DIM; i++) begin
                        updated_states[m][i] <= '0;
                        updated_cov[m][i] <= '0;
                    end
                    likelihoods[m] <= '0;
                end else if (state == ST_UPDATE_CV + m) begin
                    // Innovation (residual)
                    logic signed [STATE_WIDTH-1:0] innov [0:MEAS_DIM-1];
                    innov[0] = $signed(meas_latched[0]) - $signed(predicted_states[m][0]);
                    innov[1] = $signed(meas_latched[1]) - $signed(predicted_states[m][1]);
                    innov[2] = $signed(meas_latched[2]) - $signed(predicted_states[m][2]);
                    
                    // Innovation covariance S = H*P*H' + R (diagonal)
                    logic [STATE_WIDTH-1:0] S [0:MEAS_DIM-1];
                    S[0] = predicted_cov[m][0] + {16'b0, meas_var_latched};
                    S[1] = predicted_cov[m][1] + {16'b0, meas_var_latched};
                    S[2] = predicted_cov[m][2] + {16'b0, meas_var_latched};
                    
                    // Kalman gain K = P*H'/S (simplified for diagonal)
                    logic [STATE_WIDTH-1:0] K [0:STATE_DIM-1][0:MEAS_DIM-1];
                    for (int i = 0; i < MEAS_DIM; i++) begin
                        // K[i][i] = P[i]/S[i] for position states
                        K[i][i] = (predicted_cov[m][i] << FRAC_BITS) / S[i];
                    end
                    
                    // State update: x = x̄ + K*y
                    updated_states[m][0] <= predicted_states[m][0] + 
                        ((K[0][0] * innov[0]) >>> FRAC_BITS);
                    updated_states[m][1] <= predicted_states[m][1] + 
                        ((K[1][1] * innov[1]) >>> FRAC_BITS);
                    updated_states[m][2] <= predicted_states[m][2] + 
                        ((K[2][2] * innov[2]) >>> FRAC_BITS);
                    
                    // Velocity and acceleration: propagate from prediction
                    for (int i = 3; i < STATE_DIM; i++) begin
                        updated_states[m][i] <= predicted_states[m][i];
                    end
                    
                    // Covariance update: P = (I - K*H)*P̄
                    for (int i = 0; i < STATE_DIM; i++) begin
                        if (i < MEAS_DIM) begin
                            updated_cov[m][i] <= predicted_cov[m][i] - 
                                ((K[i][i] * predicted_cov[m][i]) >>> FRAC_BITS);
                        end else begin
                            updated_cov[m][i] <= predicted_cov[m][i];
                        end
                    end
                    
                    // Likelihood (simplified Gaussian)
                    // L = exp(-0.5 * innov' * S^-1 * innov) / sqrt(det(S))
                    logic [63:0] innov_sq_sum;
                    innov_sq_sum = (innov[0] * innov[0]) / S[0] +
                                   (innov[1] * innov[1]) / S[1] +
                                   (innov[2] * innov[2]) / S[2];
                    
                    // Approximate likelihood (higher for smaller residuals)
                    likelihoods[m] <= (32'hFFFFFFFF - innov_sq_sum[31:0]);
                end
            end
        end
    endgenerate
    
    //--------------------------------------------------------------------------
    // Model Probability Update and Output Combination
    //--------------------------------------------------------------------------
    logic [NUM_MODELS-1:0][15:0] updated_probs;
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int m = 0; m < NUM_MODELS; m++) begin
                updated_probs[m] <= 16'h5555;  // 1/3
            end
        end else if (state == ST_COMBINE) begin
            // Update probabilities: μ_j = c_j * L_j * Σ_i π_{ij} * μ_i
            // Normalize so Σ μ_j = 1
            logic [63:0] prob_sum = '0;
            logic [31:0] unnorm_probs [NUM_MODELS-1:0];
            
            for (int j = 0; j < NUM_MODELS; j++) begin
                unnorm_probs[j] = (likelihoods[j] >>> 16) * 
                    (current_track.models[j].probability);
                prob_sum = prob_sum + unnorm_probs[j];
            end
            
            // Normalize
            if (prob_sum > 0) begin
                for (int j = 0; j < NUM_MODELS; j++) begin
                    updated_probs[j] <= (unnorm_probs[j] << 16) / prob_sum[31:0];
                end
            end
            
            // Compute combined state (probability-weighted average)
            for (int s = 0; s < STATE_DIM; s++) begin
                automatic logic signed [2*STATE_WIDTH-1:0] weighted_sum = '0;
                for (int m = 0; m < NUM_MODELS; m++) begin
                    weighted_sum = weighted_sum + 
                        ($signed(updated_states[m][s]) * $signed({16'b0, updated_probs[m]}));
                end
                current_track.combined_state[s] <= weighted_sum[STATE_WIDTH+15:16];
            end
            
            // Update track models
            for (int m = 0; m < NUM_MODELS; m++) begin
                current_track.models[m].state <= updated_states[m];
                current_track.models[m].covariance <= updated_cov[m];
                current_track.models[m].probability <= updated_probs[m];
            end
        end
    end
    
    //--------------------------------------------------------------------------
    // Track Management
    //--------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int t = 0; t < MAX_TRACKS; t++) begin
                tracks[t].active <= 1'b0;
            end
        end else if (state == ST_TRACK_MGMT) begin
            // Update hit/miss counts
            current_track.hit_count <= current_track.hit_count + 1;
            
            // Confirm track if enough hits
            if (current_track.hit_count >= cfg_confirm_hits) begin
                current_track.confirmed <= 1'b1;
            end
            
            // Write back to track memory
            tracks[current_track_id] <= current_track;
        end
    end
    
    // Count active tracks
    always_comb begin
        automatic logic [5:0] count = '0;
        for (int t = 0; t < MAX_TRACKS; t++) begin
            if (tracks[t].active) count = count + 1;
        end
        num_active_tracks = count;
    end
    
    //--------------------------------------------------------------------------
    // Output
    //--------------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state_out <= '0;
            covariance_diag <= '0;
            track_id_out <= '0;
            track_valid <= 1'b0;
            model_probs <= '0;
            track_confirmed <= 1'b0;
            track_lost <= 1'b0;
        end else if (state == ST_OUTPUT) begin
            state_out <= current_track.combined_state;
            
            // Combined covariance (simplified: weighted average of diagonals)
            for (int i = 0; i < STATE_DIM; i++) begin
                automatic logic [2*STATE_WIDTH-1:0] cov_sum = '0;
                for (int m = 0; m < NUM_MODELS; m++) begin
                    cov_sum = cov_sum + (updated_cov[m][i] * updated_probs[m]);
                end
                covariance_diag[i] <= cov_sum[STATE_WIDTH+15:16];
            end
            
            track_id_out <= current_track_id;
            track_valid <= 1'b1;
            model_probs <= updated_probs;
            track_confirmed <= current_track.confirmed;
            track_lost <= 1'b0;
        end else begin
            track_valid <= 1'b0;
        end
    end
    
    //--------------------------------------------------------------------------
    // Status
    //--------------------------------------------------------------------------
    assign busy = (state != ST_IDLE);
    assign overflow = (num_active_tracks >= MAX_TRACKS);

endmodule
