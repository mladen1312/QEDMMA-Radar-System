//=============================================================================
// QEDMMA v3.2 - Multi-Bank Correlator Top (Full Range Coverage)
// [REQ-MULTIBANK-001] Instantiate N banks for extended range window
// [REQ-MULTIBANK-002] Bank tiling with configurable overlap
// [REQ-MULTIBANK-003] Unified AXI-Stream output multiplexer
//
// Author: Dr. Mladen Mešter
// Independently Validated
// Copyright (c) 2026 - All Rights Reserved
//
// Architecture:
//   Single 512-lane bank covers 384m (512 × 0.75m)
//   For tactical mode: 8 banks = 3.07 km window
//   For strategic mode: Dynamic bank allocation via range gates
//
//   ┌────────────────────────────────────────────────────────────────────┐
//   │                    MULTI-BANK CORRELATOR TOP                       │
//   ├────────────────────────────────────────────────────────────────────┤
//   │                                                                    │
//   │  ADC ──▶ Bank[0] ──▶ Lanes 0-511     (0 - 384m)                   │
//   │     └──▶ Bank[1] ──▶ Lanes 512-1023  (384m - 768m)                │
//   │     └──▶ Bank[2] ──▶ Lanes 1024-1535 (768m - 1152m)               │
//   │     └──▶ ...                                                       │
//   │     └──▶ Bank[7] ──▶ Lanes 3584-4095 (2688m - 3072m)              │
//   │                                                                    │
//   │  Optional: Range gate steering for extended range (800 km)        │
//   │                                                                    │
//   └────────────────────────────────────────────────────────────────────┘
//
// Resources (8-bank configuration):
//   LUT: ~40K (8 × 5K)
//   FF:  ~80K (8 × 10K)
//   BRAM: 0 (zero-DSP architecture)
//   DSP48: 0 (XOR-based correlation)
//
// Target: Xilinx Zynq UltraScale+ ZU47DR @ 200 MHz
//=============================================================================

`timescale 1ns / 1ps

module qedmma_correlator_bank_top #(
    parameter int NUM_BANKS       = 8,            // Number of parallel banks
    parameter int LANES_PER_BANK  = 512,          // Lanes per bank
    parameter int SAMPLE_WIDTH    = 16,           // ADC sample width
    parameter int ACC_WIDTH       = 48,           // Accumulator width
    parameter int AXI_DATA_WIDTH  = 64            // AXI-Stream width
)(
    //=========================================================================
    // Clocks and Resets
    //=========================================================================
    input  logic                          clk_fast,       // 200 MHz
    input  logic                          clk_axi,        // 100 MHz
    input  logic                          rst_n,
    
    //=========================================================================
    // ADC Input (I/Q)
    //=========================================================================
    input  logic signed [SAMPLE_WIDTH-1:0] adc_i,
    input  logic signed [SAMPLE_WIDTH-1:0] adc_q,
    input  logic                          adc_valid,
    
    //=========================================================================
    // PRBS Reference
    //=========================================================================
    input  logic                          prbs_bit,
    input  logic                          prbs_valid,
    
    //=========================================================================
    // White Rabbit Sync
    //=========================================================================
    input  logic                          wr_pps,
    input  logic                          wr_sync_enable,
    
    //=========================================================================
    // AXI-Stream Output (merged from all banks)
    //=========================================================================
    output logic [AXI_DATA_WIDTH-1:0]     m_axis_tdata,
    output logic                          m_axis_tvalid,
    output logic                          m_axis_tlast,
    output logic [3:0]                    m_axis_tid,     // Bank ID
    input  logic                          m_axis_tready,
    
    //=========================================================================
    // Configuration
    //=========================================================================
    input  logic                          cfg_enable,
    input  logic                          cfg_clear,
    input  logic [31:0]                   cfg_integration_count,
    input  logic                          cfg_dump_on_pps,
    input  logic [NUM_BANKS-1:0]          cfg_bank_enable, // Enable mask
    input  logic [31:0]                   cfg_range_gate_offset, // Extended range
    
    //=========================================================================
    // Status
    //=========================================================================
    output logic [31:0]                   status_chip_count,
    output logic [12:0]                   status_global_peak_lane, // 0-4095
    output logic [ACC_WIDTH-1:0]          status_global_peak_mag,
    output logic [2:0]                    status_peak_bank,
    output logic [NUM_BANKS-1:0]          status_bank_done,
    output logic [NUM_BANKS-1:0]          status_bank_overflow
);

    //=========================================================================
    // Local Parameters
    //=========================================================================
    localparam int TOTAL_LANES = NUM_BANKS * LANES_PER_BANK;  // 4096 for 8 banks
    localparam int LOG2_BANKS = $clog2(NUM_BANKS);
    
    //=========================================================================
    // Bank Instantiation Signals
    //=========================================================================
    
    // Per-bank AXI-Stream outputs
    logic [AXI_DATA_WIDTH-1:0] bank_tdata [NUM_BANKS];
    logic bank_tvalid [NUM_BANKS];
    logic bank_tlast [NUM_BANKS];
    logic bank_tready [NUM_BANKS];
    
    // Per-bank status
    logic [9:0] bank_peak_lane [NUM_BANKS];
    logic [ACC_WIDTH-1:0] bank_peak_mag [NUM_BANKS];
    logic bank_done [NUM_BANKS];
    logic bank_overflow [NUM_BANKS];
    
    //=========================================================================
    // Delay Line Extension for Multi-Bank
    //=========================================================================
    // Feed delayed samples to each bank for range offset
    // Bank N receives samples delayed by N × LANES_PER_BANK clocks
    
    logic signed [SAMPLE_WIDTH-1:0] bank_adc_i [NUM_BANKS];
    logic signed [SAMPLE_WIDTH-1:0] bank_adc_q [NUM_BANKS];
    logic bank_adc_valid [NUM_BANKS];
    
    // Extended delay line for bank input staging
    logic signed [SAMPLE_WIDTH-1:0] ext_delay_i [NUM_BANKS * LANES_PER_BANK];
    logic signed [SAMPLE_WIDTH-1:0] ext_delay_q [NUM_BANKS * LANES_PER_BANK];
    
    always_ff @(posedge clk_fast or negedge rst_n) begin
        if (!rst_n) begin
            for (int i = 0; i < NUM_BANKS * LANES_PER_BANK; i++) begin
                ext_delay_i[i] <= '0;
                ext_delay_q[i] <= '0;
            end
        end else if (adc_valid && cfg_enable) begin
            ext_delay_i[0] <= adc_i;
            ext_delay_q[0] <= adc_q;
            
            for (int i = 1; i < NUM_BANKS * LANES_PER_BANK; i++) begin
                ext_delay_i[i] <= ext_delay_i[i-1];
                ext_delay_q[i] <= ext_delay_q[i-1];
            end
        end
    end
    
    // Tap delay line at bank boundaries
    genvar bank;
    generate
        for (bank = 0; bank < NUM_BANKS; bank++) begin : gen_bank_taps
            localparam int TAP_OFFSET = bank * LANES_PER_BANK;
            
            assign bank_adc_i[bank] = ext_delay_i[TAP_OFFSET];
            assign bank_adc_q[bank] = ext_delay_q[TAP_OFFSET];
            assign bank_adc_valid[bank] = adc_valid && cfg_bank_enable[bank];
        end
    endgenerate
    
    //=========================================================================
    // Correlator Bank Instantiation
    //=========================================================================
    
    generate
        for (bank = 0; bank < NUM_BANKS; bank++) begin : gen_banks
            qedmma_correlator_bank_v32 #(
                .NUM_LANES(LANES_PER_BANK),
                .SAMPLE_WIDTH(SAMPLE_WIDTH),
                .ACC_WIDTH(ACC_WIDTH),
                .AXI_DATA_WIDTH(AXI_DATA_WIDTH)
            ) u_bank (
                .clk_fast(clk_fast),
                .clk_axi(clk_axi),
                .rst_n(rst_n),
                
                // ADC input (from extended delay line)
                .adc_i(bank_adc_i[bank]),
                .adc_q(bank_adc_q[bank]),
                .adc_valid(bank_adc_valid[bank]),
                
                // PRBS reference (same for all banks)
                .prbs_bit(prbs_bit),
                .prbs_valid(prbs_valid),
                
                // White Rabbit sync
                .wr_pps(wr_pps),
                .wr_sync_enable(wr_sync_enable),
                
                // AXI-Stream output
                .m_axis_tdata(bank_tdata[bank]),
                .m_axis_tvalid(bank_tvalid[bank]),
                .m_axis_tlast(bank_tlast[bank]),
                .m_axis_tready(bank_tready[bank]),
                
                // Configuration
                .cfg_enable(cfg_enable && cfg_bank_enable[bank]),
                .cfg_clear(cfg_clear),
                .cfg_integration_count(cfg_integration_count),
                .cfg_dump_on_pps(cfg_dump_on_pps),
                
                // Status
                .status_chip_count(),  // Use global counter
                .status_peak_lane(bank_peak_lane[bank]),
                .status_peak_magnitude(bank_peak_mag[bank]),
                .status_integration_done(bank_done[bank]),
                .status_overflow(bank_overflow[bank])
            );
        end
    endgenerate
    
    //=========================================================================
    // Global Peak Finder (across all banks)
    //=========================================================================
    
    logic [12:0] global_peak_lane;
    logic [ACC_WIDTH-1:0] global_peak_mag;
    logic [2:0] peak_bank_idx;
    
    always_ff @(posedge clk_fast or negedge rst_n) begin
        if (!rst_n) begin
            global_peak_lane <= '0;
            global_peak_mag <= '0;
            peak_bank_idx <= '0;
        end else begin
            // Find global maximum across all banks
            logic [ACC_WIDTH-1:0] max_mag;
            logic [2:0] max_bank;
            logic [12:0] max_lane;
            
            max_mag = bank_peak_mag[0];
            max_bank = 3'd0;
            max_lane = {3'd0, bank_peak_lane[0]};
            
            for (int b = 1; b < NUM_BANKS; b++) begin
                if (bank_peak_mag[b] > max_mag) begin
                    max_mag = bank_peak_mag[b];
                    max_bank = b[2:0];
                    max_lane = {b[2:0], bank_peak_lane[b]};
                end
            end
            
            global_peak_lane <= max_lane;
            global_peak_mag <= max_mag;
            peak_bank_idx <= max_bank;
        end
    end
    
    assign status_global_peak_lane = global_peak_lane;
    assign status_global_peak_mag = global_peak_mag;
    assign status_peak_bank = peak_bank_idx;
    
    //=========================================================================
    // AXI-Stream Output Multiplexer
    //=========================================================================
    // Round-robin arbitration across banks
    
    logic [2:0] arb_bank;
    logic arb_valid;
    
    typedef enum logic [1:0] {
        ARB_IDLE,
        ARB_TRANSMIT,
        ARB_NEXT
    } arb_state_t;
    
    arb_state_t arb_state;
    
    always_ff @(posedge clk_axi or negedge rst_n) begin
        if (!rst_n) begin
            arb_state <= ARB_IDLE;
            arb_bank <= '0;
            m_axis_tvalid <= 1'b0;
            m_axis_tlast <= 1'b0;
            m_axis_tdata <= '0;
            m_axis_tid <= '0;
        end else begin
            case (arb_state)
                ARB_IDLE: begin
                    // Find next bank with valid data
                    for (int b = 0; b < NUM_BANKS; b++) begin
                        int idx;
                        idx = (arb_bank + b) % NUM_BANKS;
                        if (bank_tvalid[idx]) begin
                            arb_bank <= idx[2:0];
                            arb_state <= ARB_TRANSMIT;
                            break;
                        end
                    end
                    m_axis_tvalid <= 1'b0;
                end
                
                ARB_TRANSMIT: begin
                    if (bank_tvalid[arb_bank]) begin
                        m_axis_tdata <= bank_tdata[arb_bank];
                        m_axis_tvalid <= 1'b1;
                        m_axis_tlast <= bank_tlast[arb_bank];
                        m_axis_tid <= arb_bank;
                        bank_tready[arb_bank] <= m_axis_tready;
                        
                        if (bank_tlast[arb_bank] && m_axis_tready) begin
                            arb_state <= ARB_NEXT;
                        end
                    end else begin
                        arb_state <= ARB_IDLE;
                    end
                end
                
                ARB_NEXT: begin
                    m_axis_tvalid <= 1'b0;
                    m_axis_tlast <= 1'b0;
                    arb_bank <= (arb_bank + 1) % NUM_BANKS;
                    arb_state <= ARB_IDLE;
                end
                
                default: arb_state <= ARB_IDLE;
            endcase
        end
    end
    
    //=========================================================================
    // Status Aggregation
    //=========================================================================
    
    // Global chip counter (from first enabled bank)
    assign status_chip_count = cfg_bank_enable[0] ? 
        gen_banks[0].u_bank.status_chip_count : '0;
    
    // Bank status aggregation
    always_comb begin
        for (int b = 0; b < NUM_BANKS; b++) begin
            status_bank_done[b] = bank_done[b];
            status_bank_overflow[b] = bank_overflow[b];
        end
    end

endmodule
